library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity conv_img_buffer is
	Port ( 
		clk : in  STD_LOGIC
	);
end conv_img_buffer;

architecture Behavioral of conv_img_buffer is

begin


end Behavioral;

