library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
library ieee_proposed;
use ieee_proposed.fixed_float_types.all;
use ieee_proposed.fixed_pkg.all;

entity convolution is
    Port ( pixel_in : in  STD_LOGIC;
           pixel_out : out  STD_LOGIC);
end convolution;

architecture Behavioral of convolution is

begin


end Behavioral;

