--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 


library IEEE;
use IEEE.STD_LOGIC_1164.all;

package custom_type_pkg is

type bit_array is array(integer range <>) of std_logic;

end custom_type_pkg;


package body custom_type_pkg is

end custom_type_pkg;
